library verilog;
use verilog.vl_types.all;
entity testbench_alterado is
end testbench_alterado;
