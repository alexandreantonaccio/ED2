library verilog;
use verilog.vl_types.all;
entity tb_relogio is
end tb_relogio;
