library verilog;
use verilog.vl_types.all;
entity relogio_tb is
end relogio_tb;
