module tb_relogio();

    // inputs
    reg reset;
    reg clk;
    reg [1:0] H_in1;
    reg [3:0] H_in0;
    reg [3:0] M_in1;
    reg [3:0] M_in0;
    reg LD_time;

    // saida do relogio principal
    wire [1:0] H_out1;
    wire [3:0] H_out0;
    wire [3:0] M_out1;
    wire [3:0] M_out0;
    wire [3:0] S_out1;
    wire [3:0] S_out0;

    // saida alternada
    wire [1:0] alt_H_out1;
    wire [3:0] alt_H_out0;
    wire [3:0] alt_M_out1;
    wire [3:0] alt_M_out0;
    wire [3:0] alt_S_out1;
    wire [3:0] alt_S_out0;

    // teste
    relogio teste (
        .reset(reset), 
        .clk(clk), 
        .H_in1(H_in1), 
        .H_in0(H_in0), 
        .M_in1(M_in1), 
        .M_in0(M_in0), 
        .LD_time(LD_time), 
        .H_out1(H_out1), 
        .H_out0(H_out0), 
        .M_out1(M_out1), 
        .M_out0(M_out0), 
        .S_out1(S_out1), 
        .S_out0(S_out0), 
        .alt_H_out1(alt_H_out1), 
        .alt_H_out0(alt_H_out0), 
        .alt_M_out1(alt_M_out1), 
        .alt_M_out0(alt_M_out0), 
        .alt_S_out1(alt_S_out1), 
        .alt_S_out0(alt_S_out0)
    );

    // gera clock
    initial begin
        clk = 0;
        forever #50000000 clk = ~clk;  // pulso 1 seg
    end

    // testa sequencia
    initial begin
        // inicializa 
        reset = 1;
        H_in1 = 1;
        H_in0 = 0;
        M_in1 = 1;
        M_in0 = 9;
        LD_time = 0;

        // reset = 0 apos 1 seg
        #100000000;
        reset = 0;

        #100000000;
        H_in1 = 1;
        H_in0 = 0;
        M_in1 = 2;
        M_in0 = 0;
        LD_time = 1;

        #100000000;
        LD_time = 0;

        repeat(86400) begin
            #1000000000;  
        end

        $stop;
    end

endmodule
