`timescale 1ns / 1ps

module relogio_tb;

    // Declara��o de sinais de entrada como reg
    reg reset;
    reg clk;
    reg [1:0] H_in1;
    reg [3:0] H_in0;
    reg [3:0] M_in1;
    reg [3:0] M_in0;
    reg LD_time;

    // Declara��o de sinais de sa�da como wire
    wire [1:0] H_out1;
    wire [3:0] H_out0;
    wire [3:0] M_out1;
    wire [3:0] M_out0;
    wire [3:0] S_out1;
    wire [3:0] S_out0;
    wire [1:0] alt_H_out1;
    wire [3:0] alt_H_out0;
    wire [3:0] alt_M_out1;
    wire [3:0] alt_M_out0;
    wire [3:0] alt_S_out1;
    wire [3:0] alt_S_out0;

    // Instancia��o do m�dulo DUT (Device Under Test)
    relogio_alterado DUT (
        .reset(reset),
        .clk(clk),
        .H_in1(H_in1),
        .H_in0(H_in0),
        .M_in1(M_in1),
        .M_in0(M_in0),
        .LD_time(LD_time),
        .H_out1(H_out1),
        .H_out0(H_out0),
        .M_out1(M_out1),
        .M_out0(M_out0),
        .S_out1(S_out1),
        .S_out0(S_out0),
        .alt_H_out1(alt_H_out1),
        .alt_H_out0(alt_H_out0),
        .alt_M_out1(alt_M_out1),
        .alt_M_out0(alt_M_out0),
        .alt_S_out1(alt_S_out1),
        .alt_S_out0(alt_S_out0)
    );

    // Gera��o do sinal de clock com per�odo de 10 ns
    initial begin
        clk = 0;
        forever #5 clk = ~clk; // Per�odo total de 10 ns
    end

    // Inicializa��o e aplica��o dos est�mulos
    initial begin
        // Inicializa��o das entradas
        reset = 1;
        H_in1 = 2'b00;   // Horas: 00
        H_in0 = 4'd0;
        M_in1 = 4'd0;    // Minutos: 00
        M_in0 = 4'd0;
        LD_time = 0;

        // Monitoramento das sa�das
        $monitor("Time=%0t | Reset=%b | LD_time=%b | H=%d%d | M=%d%d | S=%d%d | Display Mode=%b",
                 $time, reset, LD_time, H_out1, H_out0, M_out1, M_out0, S_out1, S_out0, DUT.display_modo);

        // Aplica��o do reset
        #20;
        reset = 0;

        // Carregar tempo inicial (exemplo: 12:34)
        #10;
        H_in1 = 2'b01;   // 1
        H_in0 = 4'd2;    // 2
        M_in1 = 4'd3;    // 3
        M_in0 = 4'd4;    // 4
        LD_time = 1;

        #10;
        LD_time = 0; // Desativar LD_time ap�s carregar

        // Simular a contagem de tempo
        // A quantidade de tempo simulada depender� da rela��o entre clk e clk_1s
        // Para acelerar a simula��o, voc� pode ajustar o contador interno ou os tempos de espera

        // Simula��o por um per�odo suficiente para observar a contagem
        #100000; // Tempo total de simula��o (ajuste conforme necess�rio)

        // Finaliza��o da simula��o
        $finish;
    end

    // Opcional: Dump de ondas para visualiza��o no GTKWave ou similar
    initial begin
        $dumpfile("relogio_tb.vcd");
        $dumpvars(0, relogio_tb);
    end

endmodule
