library verilog;
use verilog.vl_types.all;
entity relogio_johnson_tb is
end relogio_johnson_tb;
